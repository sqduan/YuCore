/********************************************************************************
 *                                                                              *
 *                          Yu Core - Single Cycle Version                      *
 *                                                                              *
 *------------------------------------------------------------------------------*
 * File Name   : TestParameters.vh                                              *
 * Description : This file describes the parameters of test file                *
 *               used in Yu Core                                                *
 * Author      : Shiqi Duan                                                     *
 * Date        : 2022/11/6                                                      *
*********************************************************************************/
`ifndef _TEST_PARAMETERS_VH_
`define _TEST_PARAMETERS_VH_

parameter SUCCESS = 0;

`endif